netcdf hycom1_25 {
dimensions:
	layers = 25 ;
	interfaces = 26 ;
variables:
	double dz(layers) ;
		dz:long_name = "z* coordinate level thickness" ;
		dz:units = "m" ;
	double sigma0(interfaces) ;
		sigma0:long_name = "Interface target potential density referenced to 0 dbars" ;
		sigma0:units = "kg/m3" ;
data:

 dz = 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 sigma0 = 1027, 1027.167277712, 1027.197033136, 1027.22678856, 
    1027.256543984, 1027.286299408, 1027.316054832, 1027.345810256, 
    1027.37556568, 1027.405321104, 1027.435076528, 1027.464831952, 
    1027.494587376, 1027.5243428, 1027.554098224, 1027.583853648, 
    1027.613609072, 1027.643364496, 1027.67311992, 1027.702875344, 
    1027.732630768, 1027.762386192, 1027.792141616, 1027.82189704, 
    1027.851652464, 1027.881407888 ;
}
